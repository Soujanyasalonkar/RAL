`include "seq_item.sv"
`include "reg_pkt.sv"
`include "ral_adapter.sv"

`include "base_sequence.sv"
//`include "sequencer.sv"
//`include "driver.sv"
//`include "monitor.sv"
`include "my_agent.sv"
`include "reg_env.sv"
`include "reset_seq.sv"
